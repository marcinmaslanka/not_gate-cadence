//Verilog HDL for "AMS", "not_gate" "functional"


module not_gate (y ,a );
output y;
input a;

assign y=~a;

endmodule
